`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Habib University
// Engineer: PalmPilot X Team
// 
// Create Date: 05/01/2025 05:19:22 PM
// Design Name: PalmPilot X
// Module Name: movement
// Project Name: PalmPilot X
// Target Devices: Basys 3
// Tool Versions: Vivado 2020.1
// Description: This module translates IR sensor inputs into directional text display
// 
// Dependencies: None
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Module takes 4-bit IR sensor input and displays corresponding movement text
// (FORWARD, BACKWARD, LEFT, RIGHT, combinations, or HOVER ON SENSOR)
//////////////////////////////////////////////////////////////////////////////////


module movement(
    input [3:0] ir,
    input [10:0] x,
    output reg [6:0] char_addr_TEXT
    );
    
    
    always @* begin
    char_addr_TEXT = 
    ir[0]&&ir[1]?
    (x >= 128  && x < 160)  ? 7'h49 :  // 'I'
    (x >= 160  && x < 192)  ? 7'h4E :  // 'N'
    (x >= 192  && x < 224)  ? 7'h56 :  // 'V'
    (x >= 224  && x < 256)  ? 7'h41 :  // 'A'
    (x >= 256  && x < 288)  ? 7'h4C :  // 'L'
    (x >= 288  && x < 320)  ? 7'h49 :  // 'I'
    (x >= 320  && x < 352)  ? 7'h44 :  // 'D'
    (x >= 352  && x < 384)  ? 7'h20 :  // ' '
    (x >= 384  && x < 416)  ? 7'h49 :  // 'I'
    (x >= 416  && x < 448)  ? 7'h4E :  // 'N'
    (x >= 448  && x < 480)  ? 7'h50 :  // 'P'
    (x >= 480  && x < 512)  ? 7'h55 :  // 'U'
    (x >= 512  && x < 544)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space

    :ir[2]&&ir[3]?
    (x >= 128  && x < 160)  ? 7'h49 :  // 'I'
    (x >= 160  && x < 192)  ? 7'h4E :  // 'N'
    (x >= 192  && x < 224)  ? 7'h56 :  // 'V'
    (x >= 224  && x < 256)  ? 7'h41 :  // 'A'
    (x >= 256  && x < 288)  ? 7'h4C :  // 'L'
    (x >= 288  && x < 320)  ? 7'h49 :  // 'I'
    (x >= 320  && x < 352)  ? 7'h44 :  // 'D'
    (x >= 352  && x < 384)  ? 7'h20 :  // ' '
    (x >= 384  && x < 416)  ? 7'h49 :  // 'I'
    (x >= 416  && x < 448)  ? 7'h4E :  // 'N'
    (x >= 448  && x < 480)  ? 7'h50 :  // 'P'
    (x >= 480  && x < 512)  ? 7'h55 :  // 'U'
    (x >= 512  && x < 544)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space                           
    :ir[2]&&ir[1]?
    (x >= 128  && x < 160)  ? 7'h46 :  // 'F'
    (x >= 160  && x < 192)  ? 7'h4F :  // 'O'
    (x >= 192  && x < 224)  ? 7'h52 :  // 'R'
    (x >= 224  && x < 256)  ? 7'h57 :  // 'W'
    (x >= 256  && x < 288)  ? 7'h41 :  // 'A'
    (x >= 288  && x < 320)  ? 7'h52 :  // 'R'
    (x >= 320  && x < 352)  ? 7'h44 :  // 'D'
    (x >= 352  && x < 384)  ? 7'h20 :  // ' '
    (x >= 384  && x < 416)  ? 7'h41 :  // 'A'
    (x >= 416  && x < 448)  ? 7'h4E :  // 'N'
    (x >= 448  && x < 480)  ? 7'h44 :  // 'D'
    (x >= 480  && x < 512)  ? 7'h20 :  // ' '
    (x >= 512  && x < 544)  ? 7'h52 :  // 'R'
    (x >= 544  && x < 576)  ? 7'h49 :  // 'I'
    (x >= 576  && x < 608)  ? 7'h47 :  // 'G'
    (x >= 608  && x < 640)  ? 7'h48 :  // 'H'
    (x >= 640  && x < 672)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space
    

    :ir[3]&&ir[1]?
    (x >= 128  && x < 160)  ? 7'h46 :  // 'F'
    (x >= 160  && x < 192)  ? 7'h4F :  // 'O'
    (x >= 192  && x < 224)  ? 7'h52 :  // 'R'
    (x >= 224  && x < 256)  ? 7'h57 :  // 'W'
    (x >= 256  && x < 288)  ? 7'h41 :  // 'A'
    (x >= 288  && x < 320)  ? 7'h52 :  // 'R'
    (x >= 320  && x < 352)  ? 7'h44 :  // 'D'
    (x >= 352  && x < 384)  ? 7'h20 :  // ' '
    (x >= 384  && x < 416)  ? 7'h41 :  // 'A'
    (x >= 416  && x < 448)  ? 7'h4E :  // 'N'
    (x >= 448  && x < 480)  ? 7'h44 :  // 'D'
    (x >= 480  && x < 512)  ? 7'h20 :  // ' '
    (x >= 512  && x < 544)  ? 7'h4C :  // 'L'
    (x >= 544  && x < 576)  ? 7'h45 :  // 'E'
    (x >= 576  && x < 608)  ? 7'h46 :  // 'F'
    (x >= 608  && x < 640)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space

    :ir[2]&&ir[0]?
    (x >= 128  && x < 160)  ? 7'h42 :  // 'B'
    (x >= 160  && x < 192)  ? 7'h41 :  // 'A'
    (x >= 192  && x < 224)  ? 7'h43 :  // 'C'
    (x >= 224  && x < 256)  ? 7'h4B :  // 'K'
    (x >= 256  && x < 288)  ? 7'h20 :  // ' '
    (x >= 288  && x < 320)  ? 7'h41 :  // 'A'
    (x >= 320  && x < 352)  ? 7'h4E :  // 'N'
    (x >= 352  && x < 384)  ? 7'h44 :  // 'D'
    (x >= 384  && x < 416)  ? 7'h20 :  // ' '
    (x >= 416  && x < 448)  ? 7'h52 :  // 'R'
    (x >= 448  && x < 480)  ? 7'h49 :  // 'I'
    (x >= 480  && x < 512)  ? 7'h47 :  // 'G'
    (x >= 512  && x < 544)  ? 7'h48 :  // 'H'
    (x >= 544  && x < 576)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space

    :ir[3]&&ir[0]?
    (x >= 128  && x < 160)  ? 7'h42 :  // 'B'
    (x >= 160  && x < 192)  ? 7'h41 :  // 'A'
    (x >= 192  && x < 224)  ? 7'h43 :  // 'C'
    (x >= 224  && x < 256)  ? 7'h4B :  // 'K'
    (x >= 256  && x < 288)  ? 7'h20 :  // ' '
    (x >= 288  && x < 320)  ? 7'h41 :  // 'A'
    (x >= 320  && x < 352)  ? 7'h4E :  // 'N'
    (x >= 352  && x < 384)  ? 7'h44 :  // 'D'
    (x >= 384  && x < 416)  ? 7'h20 :  // ' '
    (x >= 416  && x < 448)  ? 7'h4C :  // 'L'
    (x >= 448  && x < 480)  ? 7'h45 :  // 'E'
    (x >= 480  && x < 512)  ? 7'h46 :  // 'F'
    (x >= 512  && x < 544)  ? 7'h54 :  // 'T'
                              7'h20    // Default: space

    :ir[0]?
    (x >= 128 && x < 160)   ? 7'h42 :  // 'B'
    (x >= 160 && x < 192)   ? 7'h41 :  // 'A'
    (x >= 192 && x < 224)   ? 7'h43 :  // 'C'
    (x >= 224 && x < 256)   ? 7'h4B :  // 'K'
                              7'h20    // Default: space



    :ir[1]?
    (x >= 128 && x < 160)   ? 7'h46 :  // 'F'
    (x >= 160 && x < 192)   ? 7'h4F :  // 'O'
    (x >= 192 && x < 224)   ? 7'h52 :  // 'R'
    (x >= 224 && x < 256)   ? 7'h57 :  // 'W'
    (x >= 256 && x < 288)   ? 7'h41 :  // 'A'
    (x >= 288 && x < 320)   ? 7'h52 :  // 'R'
    (x >= 320 && x < 352)   ? 7'h44 :  // 'D'
                              7'h20    // Default: space

    :ir[2]?
    (x >= 128 && x < 160)   ? 7'h52 :  // 'R'
    (x >= 160 && x < 192)   ? 7'h49 :  // 'I'
    (x >= 192 && x < 224)   ? 7'h47 :  // 'G'
    (x >= 224 && x < 256)   ? 7'h48 :  // 'H'
    (x >= 256 && x < 288)   ? 7'h54 :  // 'T'
                              7'h20    // Default: space



    :ir[3]? 
    (x >= 128 && x < 160)   ? 7'h4C :  // 'L'
    (x >= 160 && x < 192)   ? 7'h45 :  // 'E'
    (x >= 192 && x < 224)   ? 7'h46 :  // 'F'
    (x >= 224 && x < 256)   ? 7'h54 :  // 'T'
                              7'h20    // Default: space



    :
    (x >= 128 && x < 160)   ? 7'h48 :  // 'H'
    (x >= 160 && x < 192)   ? 7'h4F :  // 'O'
    (x >= 192 && x < 224)   ? 7'h56 :  // 'V'
    (x >= 224 && x < 256)   ? 7'h45 :  // 'E'
    (x >= 256 && x < 288)   ? 7'h52 :  // 'R'
    (x >= 288 && x < 320)   ? 7'h20 :  // ' '
    (x >= 320 && x < 352)   ? 7'h4F :  // 'O'
    (x >= 352 && x < 384)   ? 7'h4E :  // 'N'
    (x >= 384 && x < 416)   ? 7'h20 :  // ' '
    (x >= 416 && x < 448)   ? 7'h53 :  // 'S'
    (x >= 448 && x < 480)   ? 7'h45 :  // 'E'
    (x >= 480 && x < 512)   ? 7'h4E :  // 'N'
    (x >= 512 && x < 544)   ? 7'h53 :  // 'S'
    (x >= 544 && x < 576)   ? 7'h4F :  // 'O'
    (x >= 576 && x < 608)   ? 7'h52 :  // 'R'
                              7'h20    // Default: space

;    end   
endmodule
